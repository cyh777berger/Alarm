// Alarm.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Alarm (
		input  wire        button1_export,   //   button1.export
		input  wire        button2_export,   //   button2.export
		input  wire        button3_export,   //   button3.export
		input  wire        clk_clk,          //       clk.clk
		output wire [31:0] display_export,   //   display.export
		output wire [15:0] display_2_export, // display_2.export
		output wire        lcd_16207_RS,     // lcd_16207.RS
		output wire        lcd_16207_RW,     //          .RW
		inout  wire [7:0]  lcd_16207_data,   //          .data
		output wire        lcd_16207_E,      //          .E
		output wire        ledg_export,      //      ledg.export
		output wire [1:0]  ledr_export,      //      ledr.export
		input  wire        reset_reset_n,    //     reset.reset_n
		input  wire [3:0]  sliders_export    //   sliders.export
	);

	wire  [31:0] cpu1_data_master_readdata;                                   // mm_interconnect_0:cpu1_data_master_readdata -> cpu1:d_readdata
	wire         cpu1_data_master_waitrequest;                                // mm_interconnect_0:cpu1_data_master_waitrequest -> cpu1:d_waitrequest
	wire         cpu1_data_master_debugaccess;                                // cpu1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu1_data_master_debugaccess
	wire  [19:0] cpu1_data_master_address;                                    // cpu1:d_address -> mm_interconnect_0:cpu1_data_master_address
	wire   [3:0] cpu1_data_master_byteenable;                                 // cpu1:d_byteenable -> mm_interconnect_0:cpu1_data_master_byteenable
	wire         cpu1_data_master_read;                                       // cpu1:d_read -> mm_interconnect_0:cpu1_data_master_read
	wire         cpu1_data_master_write;                                      // cpu1:d_write -> mm_interconnect_0:cpu1_data_master_write
	wire  [31:0] cpu1_data_master_writedata;                                  // cpu1:d_writedata -> mm_interconnect_0:cpu1_data_master_writedata
	wire  [31:0] cpu1_instruction_master_readdata;                            // mm_interconnect_0:cpu1_instruction_master_readdata -> cpu1:i_readdata
	wire         cpu1_instruction_master_waitrequest;                         // mm_interconnect_0:cpu1_instruction_master_waitrequest -> cpu1:i_waitrequest
	wire  [19:0] cpu1_instruction_master_address;                             // cpu1:i_address -> mm_interconnect_0:cpu1_instruction_master_address
	wire         cpu1_instruction_master_read;                                // cpu1:i_read -> mm_interconnect_0:cpu1_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_readdata;        // lcd_16207_0:readdata -> mm_interconnect_0:lcd_16207_0_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_16207_0_control_slave_address;         // mm_interconnect_0:lcd_16207_0_control_slave_address -> lcd_16207_0:address
	wire         mm_interconnect_0_lcd_16207_0_control_slave_read;            // mm_interconnect_0:lcd_16207_0_control_slave_read -> lcd_16207_0:read
	wire         mm_interconnect_0_lcd_16207_0_control_slave_begintransfer;   // mm_interconnect_0:lcd_16207_0_control_slave_begintransfer -> lcd_16207_0:begintransfer
	wire         mm_interconnect_0_lcd_16207_0_control_slave_write;           // mm_interconnect_0:lcd_16207_0_control_slave_write -> lcd_16207_0:write
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_writedata;       // mm_interconnect_0:lcd_16207_0_control_slave_writedata -> lcd_16207_0:writedata
	wire  [31:0] mm_interconnect_0_cpu1_debug_mem_slave_readdata;             // cpu1:debug_mem_slave_readdata -> mm_interconnect_0:cpu1_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu1_debug_mem_slave_waitrequest;          // cpu1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu1_debug_mem_slave_debugaccess;          // mm_interconnect_0:cpu1_debug_mem_slave_debugaccess -> cpu1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu1_debug_mem_slave_address;              // mm_interconnect_0:cpu1_debug_mem_slave_address -> cpu1:debug_mem_slave_address
	wire         mm_interconnect_0_cpu1_debug_mem_slave_read;                 // mm_interconnect_0:cpu1_debug_mem_slave_read -> cpu1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu1_debug_mem_slave_byteenable;           // mm_interconnect_0:cpu1_debug_mem_slave_byteenable -> cpu1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu1_debug_mem_slave_write;                // mm_interconnect_0:cpu1_debug_mem_slave_write -> cpu1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu1_debug_mem_slave_writedata;            // mm_interconnect_0:cpu1_debug_mem_slave_writedata -> cpu1:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                         // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                           // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                            // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                         // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                              // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                          // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                              // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                        // mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                          // ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                           // mm_interconnect_0:ledg_s1_address -> ledg:address
	wire         mm_interconnect_0_ledg_s1_write;                             // mm_interconnect_0:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                         // mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	wire         mm_interconnect_0_button1_s1_chipselect;                     // mm_interconnect_0:button1_s1_chipselect -> button1:chipselect
	wire  [31:0] mm_interconnect_0_button1_s1_readdata;                       // button1:readdata -> mm_interconnect_0:button1_s1_readdata
	wire   [1:0] mm_interconnect_0_button1_s1_address;                        // mm_interconnect_0:button1_s1_address -> button1:address
	wire         mm_interconnect_0_button1_s1_write;                          // mm_interconnect_0:button1_s1_write -> button1:write_n
	wire  [31:0] mm_interconnect_0_button1_s1_writedata;                      // mm_interconnect_0:button1_s1_writedata -> button1:writedata
	wire         mm_interconnect_0_button2_s1_chipselect;                     // mm_interconnect_0:button2_s1_chipselect -> button2:chipselect
	wire  [31:0] mm_interconnect_0_button2_s1_readdata;                       // button2:readdata -> mm_interconnect_0:button2_s1_readdata
	wire   [1:0] mm_interconnect_0_button2_s1_address;                        // mm_interconnect_0:button2_s1_address -> button2:address
	wire         mm_interconnect_0_button2_s1_write;                          // mm_interconnect_0:button2_s1_write -> button2:write_n
	wire  [31:0] mm_interconnect_0_button2_s1_writedata;                      // mm_interconnect_0:button2_s1_writedata -> button2:writedata
	wire  [31:0] mm_interconnect_0_sliders_s1_readdata;                       // sliders:readdata -> mm_interconnect_0:sliders_s1_readdata
	wire   [1:0] mm_interconnect_0_sliders_s1_address;                        // mm_interconnect_0:sliders_s1_address -> sliders:address
	wire         mm_interconnect_0_display_s1_chipselect;                     // mm_interconnect_0:display_s1_chipselect -> display:chipselect
	wire  [31:0] mm_interconnect_0_display_s1_readdata;                       // display:readdata -> mm_interconnect_0:display_s1_readdata
	wire   [1:0] mm_interconnect_0_display_s1_address;                        // mm_interconnect_0:display_s1_address -> display:address
	wire         mm_interconnect_0_display_s1_write;                          // mm_interconnect_0:display_s1_write -> display:write_n
	wire  [31:0] mm_interconnect_0_display_s1_writedata;                      // mm_interconnect_0:display_s1_writedata -> display:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_display_2_s1_chipselect;                   // mm_interconnect_0:display_2_s1_chipselect -> display_2:chipselect
	wire  [31:0] mm_interconnect_0_display_2_s1_readdata;                     // display_2:readdata -> mm_interconnect_0:display_2_s1_readdata
	wire   [1:0] mm_interconnect_0_display_2_s1_address;                      // mm_interconnect_0:display_2_s1_address -> display_2:address
	wire         mm_interconnect_0_display_2_s1_write;                        // mm_interconnect_0:display_2_s1_write -> display_2:write_n
	wire  [31:0] mm_interconnect_0_display_2_s1_writedata;                    // mm_interconnect_0:display_2_s1_writedata -> display_2:writedata
	wire         mm_interconnect_0_rom_s1_chipselect;                         // mm_interconnect_0:rom_s1_chipselect -> rom:chipselect
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;                           // rom:readdata -> mm_interconnect_0:rom_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;                        // mm_interconnect_0:rom_s1_debugaccess -> rom:debugaccess
	wire  [14:0] mm_interconnect_0_rom_s1_address;                            // mm_interconnect_0:rom_s1_address -> rom:address
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;                         // mm_interconnect_0:rom_s1_byteenable -> rom:byteenable
	wire         mm_interconnect_0_rom_s1_write;                              // mm_interconnect_0:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;                          // mm_interconnect_0:rom_s1_writedata -> rom:writedata
	wire         mm_interconnect_0_rom_s1_clken;                              // mm_interconnect_0:rom_s1_clken -> rom:clken
	wire         mm_interconnect_0_button3_s1_chipselect;                     // mm_interconnect_0:button3_s1_chipselect -> button3:chipselect
	wire  [31:0] mm_interconnect_0_button3_s1_readdata;                       // button3:readdata -> mm_interconnect_0:button3_s1_readdata
	wire   [1:0] mm_interconnect_0_button3_s1_address;                        // mm_interconnect_0:button3_s1_address -> button3:address
	wire         mm_interconnect_0_button3_s1_write;                          // mm_interconnect_0:button3_s1_write -> button3:write_n
	wire  [31:0] mm_interconnect_0_button3_s1_writedata;                      // mm_interconnect_0:button3_s1_writedata -> button3:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // button2:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // button1:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // button3:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu1_irq_irq;                                                // irq_mapper:sender_irq -> cpu1:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [button1:reset_n, button2:reset_n, button3:reset_n, cpu1:reset_n, display:reset_n, display_2:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, lcd_16207_0:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:cpu1_reset_reset_bridge_in_reset_reset, ram:reset, rom:reset, rst_translator:in_reset, sliders:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu1:reset_req, ram:reset_req, rom:reset_req, rst_translator:reset_req_in]
	wire         cpu1_debug_reset_request_reset;                              // cpu1:debug_reset_request -> rst_controller:reset_in1

	Alarm_button1 button1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_button1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button1_s1_readdata),   //                    .readdata
		.in_port    (button1_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                 //                 irq.irq
	);

	Alarm_button1 button2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_button2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button2_s1_readdata),   //                    .readdata
		.in_port    (button2_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	Alarm_button1 button3 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_button3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button3_s1_readdata),   //                    .readdata
		.in_port    (button3_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                 //                 irq.irq
	);

	Alarm_cpu1 cpu1 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu1_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu1_data_master_read),                              //                          .read
		.d_readdata                          (cpu1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu1_data_master_write),                             //                          .write
		.d_writedata                         (cpu1_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu1_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu1_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu1_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	Alarm_display display (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_display_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display_s1_readdata),   //                    .readdata
		.out_port   (display_export)                           // external_connection.export
	);

	Alarm_display_2 display_2 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_display_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display_2_s1_readdata),   //                    .readdata
		.out_port   (display_2_export)                           // external_connection.export
	);

	Alarm_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	Alarm_lcd_16207_0 lcd_16207_0 (
		.reset_n       (~rst_controller_reset_out_reset),                           //         reset.reset_n
		.clk           (clk_clk),                                                   //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_16207_0_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_16207_0_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_16207_0_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_16207_0_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_16207_0_control_slave_address),       //              .address
		.LCD_RS        (lcd_16207_RS),                                              //      external.export
		.LCD_RW        (lcd_16207_RW),                                              //              .export
		.LCD_data      (lcd_16207_data),                                            //              .export
		.LCD_E         (lcd_16207_E)                                                //              .export
	);

	Alarm_ledg ledg (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	Alarm_ledr ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	Alarm_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	Alarm_rom rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	Alarm_sliders sliders (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_sliders_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sliders_s1_readdata), //                    .readdata
		.in_port  (sliders_export)                         // external_connection.export
	);

	Alarm_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	Alarm_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	Alarm_mm_interconnect_0 mm_interconnect_0 (
		.clk_1_clk_clk                             (clk_clk),                                                     //                        clk_1_clk.clk
		.cpu1_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                              // cpu1_reset_reset_bridge_in_reset.reset
		.cpu1_data_master_address                  (cpu1_data_master_address),                                    //                 cpu1_data_master.address
		.cpu1_data_master_waitrequest              (cpu1_data_master_waitrequest),                                //                                 .waitrequest
		.cpu1_data_master_byteenable               (cpu1_data_master_byteenable),                                 //                                 .byteenable
		.cpu1_data_master_read                     (cpu1_data_master_read),                                       //                                 .read
		.cpu1_data_master_readdata                 (cpu1_data_master_readdata),                                   //                                 .readdata
		.cpu1_data_master_write                    (cpu1_data_master_write),                                      //                                 .write
		.cpu1_data_master_writedata                (cpu1_data_master_writedata),                                  //                                 .writedata
		.cpu1_data_master_debugaccess              (cpu1_data_master_debugaccess),                                //                                 .debugaccess
		.cpu1_instruction_master_address           (cpu1_instruction_master_address),                             //          cpu1_instruction_master.address
		.cpu1_instruction_master_waitrequest       (cpu1_instruction_master_waitrequest),                         //                                 .waitrequest
		.cpu1_instruction_master_read              (cpu1_instruction_master_read),                                //                                 .read
		.cpu1_instruction_master_readdata          (cpu1_instruction_master_readdata),                            //                                 .readdata
		.button1_s1_address                        (mm_interconnect_0_button1_s1_address),                        //                       button1_s1.address
		.button1_s1_write                          (mm_interconnect_0_button1_s1_write),                          //                                 .write
		.button1_s1_readdata                       (mm_interconnect_0_button1_s1_readdata),                       //                                 .readdata
		.button1_s1_writedata                      (mm_interconnect_0_button1_s1_writedata),                      //                                 .writedata
		.button1_s1_chipselect                     (mm_interconnect_0_button1_s1_chipselect),                     //                                 .chipselect
		.button2_s1_address                        (mm_interconnect_0_button2_s1_address),                        //                       button2_s1.address
		.button2_s1_write                          (mm_interconnect_0_button2_s1_write),                          //                                 .write
		.button2_s1_readdata                       (mm_interconnect_0_button2_s1_readdata),                       //                                 .readdata
		.button2_s1_writedata                      (mm_interconnect_0_button2_s1_writedata),                      //                                 .writedata
		.button2_s1_chipselect                     (mm_interconnect_0_button2_s1_chipselect),                     //                                 .chipselect
		.button3_s1_address                        (mm_interconnect_0_button3_s1_address),                        //                       button3_s1.address
		.button3_s1_write                          (mm_interconnect_0_button3_s1_write),                          //                                 .write
		.button3_s1_readdata                       (mm_interconnect_0_button3_s1_readdata),                       //                                 .readdata
		.button3_s1_writedata                      (mm_interconnect_0_button3_s1_writedata),                      //                                 .writedata
		.button3_s1_chipselect                     (mm_interconnect_0_button3_s1_chipselect),                     //                                 .chipselect
		.cpu1_debug_mem_slave_address              (mm_interconnect_0_cpu1_debug_mem_slave_address),              //             cpu1_debug_mem_slave.address
		.cpu1_debug_mem_slave_write                (mm_interconnect_0_cpu1_debug_mem_slave_write),                //                                 .write
		.cpu1_debug_mem_slave_read                 (mm_interconnect_0_cpu1_debug_mem_slave_read),                 //                                 .read
		.cpu1_debug_mem_slave_readdata             (mm_interconnect_0_cpu1_debug_mem_slave_readdata),             //                                 .readdata
		.cpu1_debug_mem_slave_writedata            (mm_interconnect_0_cpu1_debug_mem_slave_writedata),            //                                 .writedata
		.cpu1_debug_mem_slave_byteenable           (mm_interconnect_0_cpu1_debug_mem_slave_byteenable),           //                                 .byteenable
		.cpu1_debug_mem_slave_waitrequest          (mm_interconnect_0_cpu1_debug_mem_slave_waitrequest),          //                                 .waitrequest
		.cpu1_debug_mem_slave_debugaccess          (mm_interconnect_0_cpu1_debug_mem_slave_debugaccess),          //                                 .debugaccess
		.display_s1_address                        (mm_interconnect_0_display_s1_address),                        //                       display_s1.address
		.display_s1_write                          (mm_interconnect_0_display_s1_write),                          //                                 .write
		.display_s1_readdata                       (mm_interconnect_0_display_s1_readdata),                       //                                 .readdata
		.display_s1_writedata                      (mm_interconnect_0_display_s1_writedata),                      //                                 .writedata
		.display_s1_chipselect                     (mm_interconnect_0_display_s1_chipselect),                     //                                 .chipselect
		.display_2_s1_address                      (mm_interconnect_0_display_2_s1_address),                      //                     display_2_s1.address
		.display_2_s1_write                        (mm_interconnect_0_display_2_s1_write),                        //                                 .write
		.display_2_s1_readdata                     (mm_interconnect_0_display_2_s1_readdata),                     //                                 .readdata
		.display_2_s1_writedata                    (mm_interconnect_0_display_2_s1_writedata),                    //                                 .writedata
		.display_2_s1_chipselect                   (mm_interconnect_0_display_2_s1_chipselect),                   //                                 .chipselect
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //    jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                 .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                 .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                 .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                 .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                 .chipselect
		.lcd_16207_0_control_slave_address         (mm_interconnect_0_lcd_16207_0_control_slave_address),         //        lcd_16207_0_control_slave.address
		.lcd_16207_0_control_slave_write           (mm_interconnect_0_lcd_16207_0_control_slave_write),           //                                 .write
		.lcd_16207_0_control_slave_read            (mm_interconnect_0_lcd_16207_0_control_slave_read),            //                                 .read
		.lcd_16207_0_control_slave_readdata        (mm_interconnect_0_lcd_16207_0_control_slave_readdata),        //                                 .readdata
		.lcd_16207_0_control_slave_writedata       (mm_interconnect_0_lcd_16207_0_control_slave_writedata),       //                                 .writedata
		.lcd_16207_0_control_slave_begintransfer   (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer),   //                                 .begintransfer
		.ledg_s1_address                           (mm_interconnect_0_ledg_s1_address),                           //                          ledg_s1.address
		.ledg_s1_write                             (mm_interconnect_0_ledg_s1_write),                             //                                 .write
		.ledg_s1_readdata                          (mm_interconnect_0_ledg_s1_readdata),                          //                                 .readdata
		.ledg_s1_writedata                         (mm_interconnect_0_ledg_s1_writedata),                         //                                 .writedata
		.ledg_s1_chipselect                        (mm_interconnect_0_ledg_s1_chipselect),                        //                                 .chipselect
		.ledr_s1_address                           (mm_interconnect_0_ledr_s1_address),                           //                          ledr_s1.address
		.ledr_s1_write                             (mm_interconnect_0_ledr_s1_write),                             //                                 .write
		.ledr_s1_readdata                          (mm_interconnect_0_ledr_s1_readdata),                          //                                 .readdata
		.ledr_s1_writedata                         (mm_interconnect_0_ledr_s1_writedata),                         //                                 .writedata
		.ledr_s1_chipselect                        (mm_interconnect_0_ledr_s1_chipselect),                        //                                 .chipselect
		.ram_s1_address                            (mm_interconnect_0_ram_s1_address),                            //                           ram_s1.address
		.ram_s1_write                              (mm_interconnect_0_ram_s1_write),                              //                                 .write
		.ram_s1_readdata                           (mm_interconnect_0_ram_s1_readdata),                           //                                 .readdata
		.ram_s1_writedata                          (mm_interconnect_0_ram_s1_writedata),                          //                                 .writedata
		.ram_s1_byteenable                         (mm_interconnect_0_ram_s1_byteenable),                         //                                 .byteenable
		.ram_s1_chipselect                         (mm_interconnect_0_ram_s1_chipselect),                         //                                 .chipselect
		.ram_s1_clken                              (mm_interconnect_0_ram_s1_clken),                              //                                 .clken
		.rom_s1_address                            (mm_interconnect_0_rom_s1_address),                            //                           rom_s1.address
		.rom_s1_write                              (mm_interconnect_0_rom_s1_write),                              //                                 .write
		.rom_s1_readdata                           (mm_interconnect_0_rom_s1_readdata),                           //                                 .readdata
		.rom_s1_writedata                          (mm_interconnect_0_rom_s1_writedata),                          //                                 .writedata
		.rom_s1_byteenable                         (mm_interconnect_0_rom_s1_byteenable),                         //                                 .byteenable
		.rom_s1_chipselect                         (mm_interconnect_0_rom_s1_chipselect),                         //                                 .chipselect
		.rom_s1_clken                              (mm_interconnect_0_rom_s1_clken),                              //                                 .clken
		.rom_s1_debugaccess                        (mm_interconnect_0_rom_s1_debugaccess),                        //                                 .debugaccess
		.sliders_s1_address                        (mm_interconnect_0_sliders_s1_address),                        //                       sliders_s1.address
		.sliders_s1_readdata                       (mm_interconnect_0_sliders_s1_readdata),                       //                                 .readdata
		.sysid_qsys_0_control_slave_address        (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //       sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata       (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                 .readdata
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                       timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                 .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                 .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                 .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect)                      //                                 .chipselect
	);

	Alarm_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu1_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
